'include latch1.v'
'include latch2.v'
'include latch3.v'
'include latch4.v'
'include hazardUnit.v'
'include alu.v'
'include memory.v'
'include mux2.v'
'include mux3.v'
'include  mux4.v'
'include registerFile.v'
module top();

reg clk;
